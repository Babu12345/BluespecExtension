package myPackage;

    
    
    interface a;

    endinterface

    module mkA();
        rule RuleName(Cond);

        endrule

    endmodule
    module mkModule(InterfaceName);

    endmodule : mkModule

    typedef enum
    tagged union

endpackage